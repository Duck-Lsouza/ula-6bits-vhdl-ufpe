arithmetic_unit