comparadores