library ieee;
use ieee.std_logic_1164.all;

entity seg7_ab is
port(
    entrada  : in  std_logic_vector(5 downto 0);
    sinal    : out std_logic;                   
    saida0   : out std_logic_vector(6 downto 0);
    saida1   : out std_logic_vector(6 downto 0) 
);
end seg7_ab;

architecture arq_seg7_ab of seg7_ab is
begin

sinal <= entrada(5);

with entrada select
saida0 <=
    "1000000" when "000000",
    "1000000" when "000001", 
    "1000000" when "000010", 
    "1000000" when "000011", 
    "1000000" when "000100", 
    "1000000" when "000101", 
    "1000000" when "000110", 
    "1000000" when "000111", 
    "1000000" when "001000", 
    "1000000" when "001001", 
    "1111001" when "001010",  
    "1111001" when "001011",
    "1111001" when "001100", 
    "1111001" when "001101", 
    "1111001" when "001110", 
    "1111001" when "001111", 
    "1111001" when "010000", 
    "1111001" when "010001", 
    "1111001" when "010010", 
    "1111001" when "010011", 
    "0100100" when "010100", 
    "0100100" when "010101",
    "0100100" when "010110", 
    "0100100" when "010111", 
    "0100100" when "011000", 
    "0100100" when "011001",
    "0100100" when "011010", 
    "0100100" when "011011",
    "0100100" when "011100", 
    "0100100" when "011101", 
    "0110000" when "011110",
    "0110000" when "011111",
    "0110000" when "100000",
    "0110000" when "100001",
    "0110000" when "100010",
    "0100100" when "100011",
    "0100100" when "100100",
    "0100100" when "100101",
    "0100100" when "100110",
    "0100100" when "100111",
    "0100100" when "101000",
    "0100100" when "101001",
    "0100100" when "101010",
    "0100100" when "101011",
    "0100100" when "101100",
    "1111001" when "101101",
    "1111001" when "101110",
    "1111001" when "101111",
    "1111001" when "110000",
    "1111001" when "110001",
    "1111001" when "110010",
    "1111001" when "110011",
    "1111001" when "110100",
    "1111001" when "110101",
    "1111001" when "110110",
    "1000000" when "110111",
    "1000000" when "111000",
    "1000000" when "111001",
    "1000000" when "111010",
    "1000000" when "111011",
    "1000000" when "111100",
    "1000000" when "111101",
    "1000000" when "111110",
    "1000000" when others;  

with entrada select
saida1 <=
    "1000000" when "000000",
    "1111001" when "000001",
    "0100100" when "000010",
    "0110000" when "000011",
    "0011001" when "000100",
    "0010010" when "000101",
    "0000010" when "000110",
    "1111000" when "000111",
    "0000000" when "001000",
    "0010000" when "001001",
    "1000000" when "001010",
    "1111001" when "001011",
    "0100100" when "001100",
    "0110000" when "001101",
    "0011001" when "001110",
    "0010010" when "001111",
    "0000010" when "010000",
    "1111000" when "010001",
    "0000000" when "010010",
    "0010000" when "010011",
    "1000000" when "010100",
    "1111001" when "010101",
    "0100100" when "010110",
    "0110000" when "010111",
    "0011001" when "011000",
    "0010010" when "011001",
    "0000010" when "011010",
    "1111000" when "011011",
    "0000000" when "011100",
    "0010000" when "011101",
    "1000000" when "011110",
    "1111001" when "011111",
    "0100100" when "100000",
    "1111001" when "100001",
    "1000000" when "100010",
    "0010000" when "100011",
    "0000000" when "100100",
    "1111000" when "100101",
    "0000010" when "100110",
    "0010010" when "100111",
    "0011001" when "101000",
    "0110000" when "101001",
    "0100100" when "101010",
    "1111001" when "101011",
    "1000000" when "101100",
    "0010000" when "101101",
    "0000000" when "101110",
    "1111000" when "101111",
    "0000010" when "110000",
    "0010010" when "110001",
    "0011001" when "110010",
    "0110000" when "110011",
    "0100100" when "110100",
    "1111001" when "110101",
    "1000000" when "110110",
    "0010000" when "110111",
    "0000000" when "111000",
    "1111000" when "111001",
    "0000010" when "111010",
    "0010010" when "111011",
    "0011001" when "111100",
    "0110000" when "111101",
    "0100100" when "111110",
    "1111001" when others;   

end arq_seg7_ab;