mux_16to1