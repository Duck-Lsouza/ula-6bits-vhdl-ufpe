logic_unity