 where select